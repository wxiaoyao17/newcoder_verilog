`timescale 1ns/1ns

/* 
    VL1 四选一多路器
*/

module mux4_1(
input [1:0]d1,d2,d3,d0,
input [1:0]sel,
output[1:0]mux_out
);
//*************code***********//

//*************code***********//
endmodule