`timescale 1ns/1ns

/* 
    VL2 异步复位的串联 T 触发器
*/

module Tff_2 (
input wire data, clk, rst,
output reg q  
);
//*************code***********//


//*************code***********//
endmodule